module key_shift();
	localparam SH_NUM = 1;
	localparam SIZE = 32;

	input i_clk, i_rst; 
	input [SIZE - 1 : 0] k;


	output  
endmodule 