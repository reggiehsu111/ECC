module key_shift();
	localparam SH_NUM = 1;
	localparam SIZE = 

	input i_clk, i_rst;
	input k;

	output 
endmodule 