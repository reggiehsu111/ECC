module Top(i_rst, i_clk, a, prime, Px, Py, k, kP);
    input i_rst;
    input i_clk;
    input [3:0] a;
    input [3:0] prime;
    input [3:0] Px;
    input [3:0] Py;
    input [3:0] k;
    
    output [3:0] kP;

endmodule